* NGSPICE file created from cs_vthref_3ho.ext - technology: gf180mcuC

.subckt cs_vthref_3ho vss vdd vb
X0 a_n1460_n1696 vb vdd vdd pfet_03v3 ad=1.456p pd=6.12u as=1.456p ps=6.12u w=5.6u l=0.56u
X1 a_n2190_n6364 a_2342_n6764 vss ppolyf_u r_width=0.8u r_length=22u
X2 vdd vb a_n1460_n1696 vdd pfet_03v3 ad=1.456p pd=6.12u as=1.456p ps=6.12u w=5.6u l=0.56u
X3 vb vb vdd vdd pfet_03v3 ad=1.456p pd=6.12u as=3.64p ps=12.5u w=5.6u l=0.56u
X4 vdd vb vb vdd pfet_03v3 ad=3.64p pd=12.5u as=1.456p ps=6.12u w=5.6u l=0.56u
X5 a_n1460_n1696 vb vdd vdd pfet_03v3 ad=1.456p pd=6.12u as=3.64p ps=12.5u w=5.6u l=0.56u
X6 vdd vb vb vdd pfet_03v3 ad=1.456p pd=6.12u as=1.456p ps=6.12u w=5.6u l=0.56u
X7 vdd vb a_n1460_n1696 vdd pfet_03v3 ad=1.456p pd=6.12u as=1.456p ps=6.12u w=5.6u l=0.56u
X8 a_n2190_n6364 vss vss ppolyf_u r_width=0.8u r_length=22u
X9 vb vb vdd vdd pfet_03v3 ad=1.456p pd=6.12u as=1.456p ps=6.12u w=5.6u l=0.56u
X10 vss vss a_n1460_n1696 vss nfet_03v3 ad=3.416p pd=12.42u as=1.456p ps=6.12u w=5.6u l=0.56u
X11 vdd vb vb vdd pfet_03v3 ad=1.456p pd=6.12u as=1.456p ps=6.12u w=5.6u l=0.56u
X12 vdd vb vb vdd pfet_03v3 ad=1.456p pd=6.12u as=1.456p ps=6.12u w=5.6u l=0.56u
X13 vdd vb a_n1460_n1696 vdd pfet_03v3 ad=1.456p pd=6.12u as=1.456p ps=6.12u w=5.6u l=0.56u
X14 vss a_n1460_n1696 vb vss nfet_03v3 ad=3.416p pd=12.42u as=1.456p ps=6.12u w=5.6u l=0.56u
X15 a_n1460_n1696 vb vdd vdd pfet_03v3 ad=1.456p pd=6.12u as=1.456p ps=6.12u w=5.6u l=0.56u
X16 a_n1460_n1696 vss vss vss nfet_03v3 ad=1.456p pd=6.12u as=3.416p ps=12.42u w=5.6u l=0.56u
X17 a_n2190_n7164 vss vss ppolyf_u r_width=0.8u r_length=22u
X18 vb a_n1460_n1696 vss vss nfet_03v3 ad=1.456p pd=6.12u as=3.416p ps=12.42u w=5.6u l=0.56u
X19 vdd vb a_n1460_n1696 vdd pfet_03v3 ad=3.64p pd=12.5u as=1.456p ps=6.12u w=5.6u l=0.56u
X20 vb vb vdd vdd pfet_03v3 ad=1.456p pd=6.12u as=1.456p ps=6.12u w=5.6u l=0.56u
X21 vb vb vdd vdd pfet_03v3 ad=1.456p pd=6.12u as=1.456p ps=6.12u w=5.6u l=0.56u
X22 a_n1460_n1696 vb vdd vdd pfet_03v3 ad=1.456p pd=6.12u as=1.456p ps=6.12u w=5.6u l=0.56u
X23 a_n2190_n7164 a_2342_n6764 vss ppolyf_u r_width=0.8u r_length=22u
C0 vdd a_n2190_n7164 0.009255f
C1 vdd a_n1460_n1696 4.17843f
C2 a_n2190_n6364 a_n2190_n7164 0.017628f
C3 vdd a_2342_n6764 0.005615f
C4 vdd a_n2190_n6364 0.00389f
C5 a_n1460_n1696 vb 1.87689f
C6 vdd vb 8.342509f
C7 vb vss 5.79116f
C8 vdd vss 83.236496f
C9 a_n2190_n7164 vss 0.674688f
C10 a_2342_n6764 vss 0.682369f
C11 a_n2190_n6364 vss 0.669913f
C12 a_n1460_n1696 vss 4.73552f
.ends

